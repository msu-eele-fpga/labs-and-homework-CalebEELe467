library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.assert_pkg.all;
use work.print_pkg.all;
use work.tb_pkg.all;

entity async_conditioner is
end entity async_conditioner;

architecture async_conditioner_arch of async_conditioner is


end architecture async_conditioner_arch;